module mux_8x1_nbit 
#(parameter N=3)
(
input [N-1:0] w0, 
input [N-1:0] w1, 
input [N-1:0] w2, 
input [N-1:0] w3, 
input [N-1:0] w4, 
input [N-1:0] w5, 
input [N-1:0] w6, 
input [N-1:0] w7, 
input [2:0] s, 
output reg [N-1:0] f
); 

always@(*)
begin




end
endmodule